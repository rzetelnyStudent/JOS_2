`define LD   3'b001  // Load: B
`define ADD  3'b010  // Add: sum of A, B and carry
`define SUB  3'b011  // Subtract: A minus B and borrow
`define NOT  3'b100  // Not: bitwise negation of A
`define AND  3'b101  // And: bitwise AND of A and B
`define OR   3'b110  // Or: bitwise OR of A and B
`define XOR  3'b111  // Xor: bitwise XOR of A and B