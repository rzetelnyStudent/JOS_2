class scoreboard;

function new();
endfunction

endclass